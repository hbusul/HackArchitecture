library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Ram512_tb is
end entity Ram512_tb;

architecture RTL of Ram512_tb is
	signal s_clk    : std_logic;
	signal s_output : std_logic_vector(15 downto 0);
	signal s_load   : std_logic := '0';
	signal s_input  : std_logic_vector(15 downto 0);
	signal s_finished : std_logic := '0';
	signal s_address : std_logic_vector(8 downto 0);
	
	type pattern_type is record
		input : std_logic_vector(15 downto 0);
		load : std_logic;
		address : std_logic_vector(8 downto 0);
		output : std_logic_vector(15 downto 0);
	end record;
	
	type pattern_array is array (natural range <>) of pattern_type;
	
	
begin
	clock_inst : entity work.ClockGenerator
		generic map(PERIOD => 20 ns)
		port map(finished => s_finished,
		clk => s_clk);
		
		RAM512: entity work.Ram512
		port map(
			clk     => s_clk,
			rst     => '0',
			load    => s_load,
			address => s_address,
			input   => s_input,
			output  => s_output
		);
	
	process
		constant patterns : pattern_array := (
			("0000000000000000",'0',"000000000","0000000000000000"),
			("0000000000000000",'0',"000000000","0000000000000000"),
			("0000000000000000",'1',"000000000","0000000000000000"),
			("0000000000000000",'1',"000000000","0000000000000000"),
			("0011001100101011",'0',"000000000","0000000000000000"),
			("0011001100101011",'0',"000000000","0000000000000000"),
			("0011001100101011",'1',"010000010","0000000000000000"),
			("0011001100101011",'1',"010000010","0011001100101011"),
			("0011001100101011",'0',"000000000","0000000000000000"),
			("0011001100101011",'0',"000000000","0000000000000000"),
			("0001001001111001",'0',"111011000","0000000000000000"),
			("0001001001111001",'0',"111011000","0000000000000000"),
			("0001001001111001",'1',"111011000","0000000000000000"),
			("0001001001111001",'1',"111011000","0001001001111001"),
			("0001001001111001",'0',"111011000","0001001001111001"),
			("0001001001111001",'0',"111011000","0001001001111001"),
			("0001001001111001",'0',"010000010","0011001100101011"),
			("0001001111111111",'0',"010000010","0011001100101011"),
			("0001001111111111",'0',"010000010","0011001100101011"),
			("0001001111111111",'1',"111111111","0000000000000000"),
			("0001001111111111",'1',"111111111","0001001111111111"),
			("0001001111111111",'0',"111111111","0001001111111111"),
			("0001001111111111",'0',"111111111","0001001111111111"),
			("0001001111111111",'0',"111011000","0001001001111001"),
			("0001001111111111",'0',"111111111","0001001111111111"),
			("0001001111111111",'0',"010101000","0000000000000000"),
			("0001001111111111",'0',"010101000","0000000000000000"),
			("0001001111111111",'0',"010101001","0000000000000000"),
			("0001001111111111",'0',"010101010","0000000000000000"),
			("0001001111111111",'0',"010101011","0000000000000000"),
			("0001001111111111",'0',"010101100","0000000000000000"),
			("0001001111111111",'0',"010101101","0000000000000000"),
			("0001001111111111",'0',"010101110","0000000000000000"),
			("0001001111111111",'0',"010101111","0000000000000000"),
			("0101010101010101",'1',"010101000","0000000000000000"),
			("0101010101010101",'1',"010101000","0101010101010101"),
			("0101010101010101",'1',"010101001","0000000000000000"),
			("0101010101010101",'1',"010101001","0101010101010101"),
			("0101010101010101",'1',"010101010","0000000000000000"),
			("0101010101010101",'1',"010101010","0101010101010101"),
			("0101010101010101",'1',"010101011","0000000000000000"),
			("0101010101010101",'1',"010101011","0101010101010101"),
			("0101010101010101",'1',"010101100","0000000000000000"),
			("0101010101010101",'1',"010101100","0101010101010101"),
			("0101010101010101",'1',"010101101","0000000000000000"),
			("0101010101010101",'1',"010101101","0101010101010101"),
			("0101010101010101",'1',"010101110","0000000000000000"),
			("0101010101010101",'1',"010101110","0101010101010101"),
			("0101010101010101",'1',"010101111","0000000000000000"),
			("0101010101010101",'1',"010101111","0101010101010101"),
			("0101010101010101",'0',"010101000","0101010101010101"),
			("0101010101010101",'0',"010101000","0101010101010101"),
			("0101010101010101",'0',"010101001","0101010101010101"),
			("0101010101010101",'0',"010101010","0101010101010101"),
			("0101010101010101",'0',"010101011","0101010101010101"),
			("0101010101010101",'0',"010101100","0101010101010101"),
			("0101010101010101",'0',"010101101","0101010101010101"),
			("0101010101010101",'0',"010101110","0101010101010101"),
			("0101010101010101",'0',"010101111","0101010101010101"),
			("1010101010101010",'1',"010101000","0101010101010101"),
			("1010101010101010",'1',"010101000","1010101010101010"),
			("1010101010101010",'0',"010101000","1010101010101010"),
			("1010101010101010",'0',"010101000","1010101010101010"),
			("1010101010101010",'0',"010101001","0101010101010101"),
			("1010101010101010",'0',"010101010","0101010101010101"),
			("1010101010101010",'0',"010101011","0101010101010101"),
			("1010101010101010",'0',"010101100","0101010101010101"),
			("1010101010101010",'0',"010101101","0101010101010101"),
			("1010101010101010",'0',"010101110","0101010101010101"),
			("1010101010101010",'0',"010101111","0101010101010101"),
			("0101010101010101",'1',"010101000","1010101010101010"),
			("0101010101010101",'1',"010101000","0101010101010101"),
			("1010101010101010",'1',"010101001","0101010101010101"),
			("1010101010101010",'1',"010101001","1010101010101010"),
			("1010101010101010",'0',"010101000","0101010101010101"),
			("1010101010101010",'0',"010101000","0101010101010101"),
			("1010101010101010",'0',"010101001","1010101010101010"),
			("1010101010101010",'0',"010101010","0101010101010101"),
			("1010101010101010",'0',"010101011","0101010101010101"),
			("1010101010101010",'0',"010101100","0101010101010101"),
			("1010101010101010",'0',"010101101","0101010101010101"),
			("1010101010101010",'0',"010101110","0101010101010101"),
			("1010101010101010",'0',"010101111","0101010101010101"),
			("0101010101010101",'1',"010101001","1010101010101010"),
			("0101010101010101",'1',"010101001","0101010101010101"),
			("1010101010101010",'1',"010101010","0101010101010101"),
			("1010101010101010",'1',"010101010","1010101010101010"),
			("1010101010101010",'0',"010101000","0101010101010101"),
			("1010101010101010",'0',"010101000","0101010101010101"),
			("1010101010101010",'0',"010101001","0101010101010101"),
			("1010101010101010",'0',"010101010","1010101010101010"),
			("1010101010101010",'0',"010101011","0101010101010101"),
			("1010101010101010",'0',"010101100","0101010101010101"),
			("1010101010101010",'0',"010101101","0101010101010101"),
			("1010101010101010",'0',"010101110","0101010101010101"),
			("1010101010101010",'0',"010101111","0101010101010101"),
			("0101010101010101",'1',"010101010","1010101010101010"),
			("0101010101010101",'1',"010101010","0101010101010101"),
			("1010101010101010",'1',"010101011","0101010101010101"),
			("1010101010101010",'1',"010101011","1010101010101010"),
			("1010101010101010",'0',"010101000","0101010101010101"),
			("1010101010101010",'0',"010101000","0101010101010101"),
			("1010101010101010",'0',"010101001","0101010101010101"),
			("1010101010101010",'0',"010101010","0101010101010101"),
			("1010101010101010",'0',"010101011","1010101010101010"),
			("1010101010101010",'0',"010101100","0101010101010101"),
			("1010101010101010",'0',"010101101","0101010101010101"),
			("1010101010101010",'0',"010101110","0101010101010101"),
			("1010101010101010",'0',"010101111","0101010101010101"),
			("0101010101010101",'1',"010101011","1010101010101010"),
			("0101010101010101",'1',"010101011","0101010101010101"),
			("1010101010101010",'1',"010101100","0101010101010101"),
			("1010101010101010",'1',"010101100","1010101010101010"),
			("1010101010101010",'0',"010101000","0101010101010101"),
			("1010101010101010",'0',"010101000","0101010101010101"),
			("1010101010101010",'0',"010101001","0101010101010101"),
			("1010101010101010",'0',"010101010","0101010101010101"),
			("1010101010101010",'0',"010101011","0101010101010101"),
			("1010101010101010",'0',"010101100","1010101010101010"),
			("1010101010101010",'0',"010101101","0101010101010101"),
			("1010101010101010",'0',"010101110","0101010101010101"),
			("1010101010101010",'0',"010101111","0101010101010101"),
			("0101010101010101",'1',"010101100","1010101010101010"),
			("0101010101010101",'1',"010101100","0101010101010101"),
			("1010101010101010",'1',"010101101","0101010101010101"),
			("1010101010101010",'1',"010101101","1010101010101010"),
			("1010101010101010",'0',"010101000","0101010101010101"),
			("1010101010101010",'0',"010101000","0101010101010101"),
			("1010101010101010",'0',"010101001","0101010101010101"),
			("1010101010101010",'0',"010101010","0101010101010101"),
			("1010101010101010",'0',"010101011","0101010101010101"),
			("1010101010101010",'0',"010101100","0101010101010101"),
			("1010101010101010",'0',"010101101","1010101010101010"),
			("1010101010101010",'0',"010101110","0101010101010101"),
			("1010101010101010",'0',"010101111","0101010101010101"),
			("0101010101010101",'1',"010101101","1010101010101010"),
			("0101010101010101",'1',"010101101","0101010101010101"),
			("1010101010101010",'1',"010101110","0101010101010101"),
			("1010101010101010",'1',"010101110","1010101010101010"),
			("1010101010101010",'0',"010101000","0101010101010101"),
			("1010101010101010",'0',"010101000","0101010101010101"),
			("1010101010101010",'0',"010101001","0101010101010101"),
			("1010101010101010",'0',"010101010","0101010101010101"),
			("1010101010101010",'0',"010101011","0101010101010101"),
			("1010101010101010",'0',"010101100","0101010101010101"),
			("1010101010101010",'0',"010101101","0101010101010101"),
			("1010101010101010",'0',"010101110","1010101010101010"),
			("1010101010101010",'0',"010101111","0101010101010101"),
			("0101010101010101",'1',"010101110","1010101010101010"),
			("0101010101010101",'1',"010101110","0101010101010101"),
			("1010101010101010",'1',"010101111","0101010101010101"),
			("1010101010101010",'1',"010101111","1010101010101010"),
			("1010101010101010",'0',"010101000","0101010101010101"),
			("1010101010101010",'0',"010101000","0101010101010101"),
			("1010101010101010",'0',"010101001","0101010101010101"),
			("1010101010101010",'0',"010101010","0101010101010101"),
			("1010101010101010",'0',"010101011","0101010101010101"),
			("1010101010101010",'0',"010101100","0101010101010101"),
			("1010101010101010",'0',"010101101","0101010101010101"),
			("1010101010101010",'0',"010101110","0101010101010101"),
			("1010101010101010",'0',"010101111","1010101010101010"),
			("0101010101010101",'1',"010101111","1010101010101010"),
			("0101010101010101",'1',"010101111","0101010101010101"),
			("0101010101010101",'0',"010101000","0101010101010101"),
			("0101010101010101",'0',"010101000","0101010101010101"),
			("0101010101010101",'0',"010101001","0101010101010101"),
			("0101010101010101",'0',"010101010","0101010101010101"),
			("0101010101010101",'0',"010101011","0101010101010101"),
			("0101010101010101",'0',"010101100","0101010101010101"),
			("0101010101010101",'0',"010101101","0101010101010101"),
			("0101010101010101",'0',"010101110","0101010101010101"),
			("0101010101010101",'0',"010101111","0101010101010101"),
			("0101010101010101",'0',"000101010","0000000000000000"),
			("0101010101010101",'0',"000101010","0000000000000000"),
			("0101010101010101",'0',"001101010","0000000000000000"),
			("0101010101010101",'0',"010101010","0101010101010101"),
			("0101010101010101",'0',"011101010","0000000000000000"),
			("0101010101010101",'0',"100101010","0000000000000000"),
			("0101010101010101",'0',"101101010","0000000000000000"),
			("0101010101010101",'0',"110101010","0000000000000000"),
			("0101010101010101",'0',"111101010","0000000000000000"),
			("0101010101010101",'1',"000101010","0000000000000000"),
			("0101010101010101",'1',"000101010","0101010101010101"),
			("0101010101010101",'1',"001101010","0000000000000000"),
			("0101010101010101",'1',"001101010","0101010101010101"),
			("0101010101010101",'1',"010101010","0101010101010101"),
			("0101010101010101",'1',"010101010","0101010101010101"),
			("0101010101010101",'1',"011101010","0000000000000000"),
			("0101010101010101",'1',"011101010","0101010101010101"),
			("0101010101010101",'1',"100101010","0000000000000000"),
			("0101010101010101",'1',"100101010","0101010101010101"),
			("0101010101010101",'1',"101101010","0000000000000000"),
			("0101010101010101",'1',"101101010","0101010101010101"),
			("0101010101010101",'1',"110101010","0000000000000000"),
			("0101010101010101",'1',"110101010","0101010101010101"),
			("0101010101010101",'1',"111101010","0000000000000000"),
			("0101010101010101",'1',"111101010","0101010101010101"),
			("0101010101010101",'0',"000101010","0101010101010101"),
			("0101010101010101",'0',"000101010","0101010101010101"),
			("0101010101010101",'0',"001101010","0101010101010101"),
			("0101010101010101",'0',"010101010","0101010101010101"),
			("0101010101010101",'0',"011101010","0101010101010101"),
			("0101010101010101",'0',"100101010","0101010101010101"),
			("0101010101010101",'0',"101101010","0101010101010101"),
			("0101010101010101",'0',"110101010","0101010101010101"),
			("0101010101010101",'0',"111101010","0101010101010101"),
			("1010101010101010",'1',"000101010","0101010101010101"),
			("1010101010101010",'1',"000101010","1010101010101010"),
			("1010101010101010",'0',"000101010","1010101010101010"),
			("1010101010101010",'0',"000101010","1010101010101010"),
			("1010101010101010",'0',"001101010","0101010101010101"),
			("1010101010101010",'0',"010101010","0101010101010101"),
			("1010101010101010",'0',"011101010","0101010101010101"),
			("1010101010101010",'0',"100101010","0101010101010101"),
			("1010101010101010",'0',"101101010","0101010101010101"),
			("1010101010101010",'0',"110101010","0101010101010101"),
			("1010101010101010",'0',"111101010","0101010101010101"),
			("0101010101010101",'1',"000101010","1010101010101010"),
			("0101010101010101",'1',"000101010","0101010101010101"),
			("1010101010101010",'1',"001101010","0101010101010101"),
			("1010101010101010",'1',"001101010","1010101010101010"),
			("1010101010101010",'0',"000101010","0101010101010101"),
			("1010101010101010",'0',"000101010","0101010101010101"),
			("1010101010101010",'0',"001101010","1010101010101010"),
			("1010101010101010",'0',"010101010","0101010101010101"),
			("1010101010101010",'0',"011101010","0101010101010101"),
			("1010101010101010",'0',"100101010","0101010101010101"),
			("1010101010101010",'0',"101101010","0101010101010101"),
			("1010101010101010",'0',"110101010","0101010101010101"),
			("1010101010101010",'0',"111101010","0101010101010101"),
			("0101010101010101",'1',"001101010","1010101010101010"),
			("0101010101010101",'1',"001101010","0101010101010101"),
			("1010101010101010",'1',"010101010","0101010101010101"),
			("1010101010101010",'1',"010101010","1010101010101010"),
			("1010101010101010",'0',"000101010","0101010101010101"),
			("1010101010101010",'0',"000101010","0101010101010101"),
			("1010101010101010",'0',"001101010","0101010101010101"),
			("1010101010101010",'0',"010101010","1010101010101010"),
			("1010101010101010",'0',"011101010","0101010101010101"),
			("1010101010101010",'0',"100101010","0101010101010101"),
			("1010101010101010",'0',"101101010","0101010101010101"),
			("1010101010101010",'0',"110101010","0101010101010101"),
			("1010101010101010",'0',"111101010","0101010101010101"),
			("0101010101010101",'1',"010101010","1010101010101010"),
			("0101010101010101",'1',"010101010","0101010101010101"),
			("1010101010101010",'1',"011101010","0101010101010101"),
			("1010101010101010",'1',"011101010","1010101010101010"),
			("1010101010101010",'0',"000101010","0101010101010101"),
			("1010101010101010",'0',"000101010","0101010101010101"),
			("1010101010101010",'0',"001101010","0101010101010101"),
			("1010101010101010",'0',"010101010","0101010101010101"),
			("1010101010101010",'0',"011101010","1010101010101010"),
			("1010101010101010",'0',"100101010","0101010101010101"),
			("1010101010101010",'0',"101101010","0101010101010101"),
			("1010101010101010",'0',"110101010","0101010101010101"),
			("1010101010101010",'0',"111101010","0101010101010101"),
			("0101010101010101",'1',"011101010","1010101010101010"),
			("0101010101010101",'1',"011101010","0101010101010101"),
			("1010101010101010",'1',"100101010","0101010101010101"),
			("1010101010101010",'1',"100101010","1010101010101010"),
			("1010101010101010",'0',"000101010","0101010101010101"),
			("1010101010101010",'0',"000101010","0101010101010101"),
			("1010101010101010",'0',"001101010","0101010101010101"),
			("1010101010101010",'0',"010101010","0101010101010101"),
			("1010101010101010",'0',"011101010","0101010101010101"),
			("1010101010101010",'0',"100101010","1010101010101010"),
			("1010101010101010",'0',"101101010","0101010101010101"),
			("1010101010101010",'0',"110101010","0101010101010101"),
			("1010101010101010",'0',"111101010","0101010101010101"),
			("0101010101010101",'1',"100101010","1010101010101010"),
			("0101010101010101",'1',"100101010","0101010101010101"),
			("1010101010101010",'1',"101101010","0101010101010101"),
			("1010101010101010",'1',"101101010","1010101010101010"),
			("1010101010101010",'0',"000101010","0101010101010101"),
			("1010101010101010",'0',"000101010","0101010101010101"),
			("1010101010101010",'0',"001101010","0101010101010101"),
			("1010101010101010",'0',"010101010","0101010101010101"),
			("1010101010101010",'0',"011101010","0101010101010101"),
			("1010101010101010",'0',"100101010","0101010101010101"),
			("1010101010101010",'0',"101101010","1010101010101010"),
			("1010101010101010",'0',"110101010","0101010101010101"),
			("1010101010101010",'0',"111101010","0101010101010101"),
			("0101010101010101",'1',"101101010","1010101010101010"),
			("0101010101010101",'1',"101101010","0101010101010101"),
			("1010101010101010",'1',"110101010","0101010101010101"),
			("1010101010101010",'1',"110101010","1010101010101010"),
			("1010101010101010",'0',"000101010","0101010101010101"),
			("1010101010101010",'0',"000101010","0101010101010101"),
			("1010101010101010",'0',"001101010","0101010101010101"),
			("1010101010101010",'0',"010101010","0101010101010101"),
			("1010101010101010",'0',"011101010","0101010101010101"),
			("1010101010101010",'0',"100101010","0101010101010101"),
			("1010101010101010",'0',"101101010","0101010101010101"),
			("1010101010101010",'0',"110101010","1010101010101010"),
			("1010101010101010",'0',"111101010","0101010101010101"),
			("0101010101010101",'1',"110101010","1010101010101010"),
			("0101010101010101",'1',"110101010","0101010101010101"),
			("1010101010101010",'1',"111101010","0101010101010101"),
			("1010101010101010",'1',"111101010","1010101010101010"),
			("1010101010101010",'0',"000101010","0101010101010101"),
			("1010101010101010",'0',"000101010","0101010101010101"),
			("1010101010101010",'0',"001101010","0101010101010101"),
			("1010101010101010",'0',"010101010","0101010101010101"),
			("1010101010101010",'0',"011101010","0101010101010101"),
			("1010101010101010",'0',"100101010","0101010101010101"),
			("1010101010101010",'0',"101101010","0101010101010101"),
			("1010101010101010",'0',"110101010","0101010101010101"),
			("1010101010101010",'0',"111101010","1010101010101010"),
			("0101010101010101",'1',"111101010","1010101010101010"),
			("0101010101010101",'1',"111101010","0101010101010101"),
			("0101010101010101",'0',"000101010","0101010101010101"),
			("0101010101010101",'0',"000101010","0101010101010101"),
			("0101010101010101",'0',"001101010","0101010101010101"),
			("0101010101010101",'0',"010101010","0101010101010101"),
			("0101010101010101",'0',"011101010","0101010101010101"),
			("0101010101010101",'0',"100101010","0101010101010101"),
			("0101010101010101",'0',"101101010","0101010101010101"),
			("0101010101010101",'0',"110101010","0101010101010101"),
			("0101010101010101",'0',"111101010","0101010101010101")
			);
		
	begin

		for i in patterns'range loop
			s_input <= patterns(i).input;
			s_load <= patterns(i).load;
			s_address <= patterns(i).address;
			wait for 60 ns;
			assert s_output = patterns(i).output
			report "bad output" severity error;
		end loop;
	

		assert false report "end of test" severity note;
		s_finished <= '1';	
		wait;
	
	end process;

end architecture RTL;
