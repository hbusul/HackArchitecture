library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Ram64_tb is
end entity Ram64_tb;

architecture RTL of Ram64_tb is
	signal s_clk    : std_logic;
	signal s_output : std_logic_vector(15 downto 0);
	signal s_load   : std_logic := '0';
	signal s_input  : std_logic_vector(15 downto 0);
	signal s_finished : std_logic := '0';
	signal s_address : std_logic_vector(5 downto 0);
	
	type pattern_type is record
		input : std_logic_vector(15 downto 0);
		load : std_logic;
		address : std_logic_vector(5 downto 0);
		output : std_logic_vector(15 downto 0);
	end record;
	
	type pattern_array is array (natural range <>) of pattern_type;
	
	
begin
	clock_inst : entity work.ClockGenerator
		generic map(PERIOD => 20 ns)
		port map(finished => s_finished,
		clk => s_clk);
		
		RAM64: entity work.Ram64
		port map(
			clk     => s_clk,
			rst     => '0',
			load    => s_load,
			address => s_address,
			input   => s_input,
			output  => s_output
		);
	
	process
		constant patterns : pattern_array := (
			("0000000000000000",'0',"000000","0000000000000000"),
			("0000000000000000",'1',"000000","0000000000000000"),
			("0000000000000000",'1',"000000","0000000000000000"),
			("0000000000000000",'1',"000000","0000000000000000"),
			("0000010100100001",'0',"000000","0000000000000000"),
			("0000010100100001",'0',"000000","0000000000000000"),
			("0000010100100001",'1',"001101","0000000000000000"),
			("0000010100100001",'1',"001101","0000010100100001"),
			("0000010100100001",'0',"000000","0000000000000000"),
			("0000010100100001",'0',"000000","0000000000000000"),
			("0001001010001011",'0',"101111","0000000000000000"),
			("0001001010001011",'0',"101111","0000000000000000"),
			("0001001010001011",'1',"101111","0000000000000000"),
			("0001001010001011",'1',"101111","0001001010001011"),
			("0001001010001011",'0',"101111","0001001010001011"),
			("0001001010001011",'0',"101111","0001001010001011"),
			("0001001010001011",'0',"001101","0000010100100001"),
			("0001100011011011",'0',"001101","0000010100100001"),
			("0001100011011011",'0',"001101","0000010100100001"),
			("0001100011011011",'1',"111111","0000000000000000"),
			("0001100011011011",'1',"111111","0001100011011011"),
			("0001100011011011",'0',"111111","0001100011011011"),
			("0001100011011011",'0',"111111","0001100011011011"),
			("0001100011011011",'0',"101111","0001001010001011"),
			("0001100011011011",'0',"111111","0001100011011011"),
			("0001100011011011",'0',"101000","0000000000000000"),
			("0001100011011011",'0',"101000","0000000000000000"),
			("0001100011011011",'0',"101001","0000000000000000"),
			("0001100011011011",'0',"101010","0000000000000000"),
			("0001100011011011",'0',"101011","0000000000000000"),
			("0001100011011011",'0',"101100","0000000000000000"),
			("0001100011011011",'0',"101101","0000000000000000"),
			("0001100011011011",'0',"101110","0000000000000000"),
			("0001100011011011",'0',"101111","0001001010001011"),
			("0101010101010101",'1',"101000","0000000000000000"),
			("0101010101010101",'1',"101000","0101010101010101"),
			("0101010101010101",'1',"101001","0000000000000000"),
			("0101010101010101",'1',"101001","0101010101010101"),
			("0101010101010101",'1',"101010","0000000000000000"),
			("0101010101010101",'1',"101010","0101010101010101"),
			("0101010101010101",'1',"101011","0000000000000000"),
			("0101010101010101",'1',"101011","0101010101010101"),
			("0101010101010101",'1',"101100","0000000000000000"),
			("0101010101010101",'1',"101100","0101010101010101"),
			("0101010101010101",'1',"101101","0000000000000000"),
			("0101010101010101",'1',"101101","0101010101010101"),
			("0101010101010101",'1',"101110","0000000000000000"),
			("0101010101010101",'1',"101110","0101010101010101"),
			("0101010101010101",'1',"101111","0001001010001011"),
			("0101010101010101",'1',"101111","0101010101010101"),
			("0101010101010101",'0',"101000","0101010101010101"),
			("0101010101010101",'0',"101000","0101010101010101"),
			("0101010101010101",'0',"101001","0101010101010101"),
			("0101010101010101",'0',"101010","0101010101010101"),
			("0101010101010101",'0',"101011","0101010101010101"),
			("0101010101010101",'0',"101100","0101010101010101"),
			("0101010101010101",'0',"101101","0101010101010101"),
			("0101010101010101",'0',"101110","0101010101010101"),
			("0101010101010101",'0',"101111","0101010101010101"),
			("1010101010101010",'1',"101000","0101010101010101"),
			("1010101010101010",'1',"101000","1010101010101010"),
			("1010101010101010",'0',"101000","1010101010101010"),
			("1010101010101010",'0',"101000","1010101010101010"),
			("1010101010101010",'0',"101001","0101010101010101"),
			("1010101010101010",'0',"101010","0101010101010101"),
			("1010101010101010",'0',"101011","0101010101010101"),
			("1010101010101010",'0',"101100","0101010101010101"),
			("1010101010101010",'0',"101101","0101010101010101"),
			("1010101010101010",'0',"101110","0101010101010101"),
			("1010101010101010",'0',"101111","0101010101010101"),
			("0101010101010101",'1',"101000","1010101010101010"),
			("0101010101010101",'1',"101000","0101010101010101"),
			("1010101010101010",'1',"101001","0101010101010101"),
			("1010101010101010",'1',"101001","1010101010101010"),
			("1010101010101010",'0',"101000","0101010101010101"),
			("1010101010101010",'0',"101000","0101010101010101"),
			("1010101010101010",'0',"101001","1010101010101010"),
			("1010101010101010",'0',"101010","0101010101010101"),
			("1010101010101010",'0',"101011","0101010101010101"),
			("1010101010101010",'0',"101100","0101010101010101"),
			("1010101010101010",'0',"101101","0101010101010101"),
			("1010101010101010",'0',"101110","0101010101010101"),
			("1010101010101010",'0',"101111","0101010101010101"),
			("0101010101010101",'1',"101001","1010101010101010"),
			("0101010101010101",'1',"101001","0101010101010101"),
			("1010101010101010",'1',"101010","0101010101010101"),
			("1010101010101010",'1',"101010","1010101010101010"),
			("1010101010101010",'0',"101000","0101010101010101"),
			("1010101010101010",'0',"101000","0101010101010101"),
			("1010101010101010",'0',"101001","0101010101010101"),
			("1010101010101010",'0',"101010","1010101010101010"),
			("1010101010101010",'0',"101011","0101010101010101"),
			("1010101010101010",'0',"101100","0101010101010101"),
			("1010101010101010",'0',"101101","0101010101010101"),
			("1010101010101010",'0',"101110","0101010101010101"),
			("1010101010101010",'0',"101111","0101010101010101"),
			("0101010101010101",'1',"101010","1010101010101010"),
			("0101010101010101",'1',"101010","0101010101010101"),
			("1010101010101010",'1',"101011","0101010101010101"),
			("1010101010101010",'1',"101011","1010101010101010"),
			("1010101010101010",'0',"101000","0101010101010101"),
			("1010101010101010",'0',"101000","0101010101010101"),
			("1010101010101010",'0',"101001","0101010101010101"),
			("1010101010101010",'0',"101010","0101010101010101"),
			("1010101010101010",'0',"101011","1010101010101010"),
			("1010101010101010",'0',"101100","0101010101010101"),
			("1010101010101010",'0',"101101","0101010101010101"),
			("1010101010101010",'0',"101110","0101010101010101"),
			("1010101010101010",'0',"101111","0101010101010101"),
			("0101010101010101",'1',"101011","1010101010101010"),
			("0101010101010101",'1',"101011","0101010101010101"),
			("1010101010101010",'1',"101100","0101010101010101"),
			("1010101010101010",'1',"101100","1010101010101010"),
			("1010101010101010",'0',"101000","0101010101010101"),
			("1010101010101010",'0',"101000","0101010101010101"),
			("1010101010101010",'0',"101001","0101010101010101"),
			("1010101010101010",'0',"101010","0101010101010101"),
			("1010101010101010",'0',"101011","0101010101010101"),
			("1010101010101010",'0',"101100","1010101010101010"),
			("1010101010101010",'0',"101101","0101010101010101"),
			("1010101010101010",'0',"101110","0101010101010101"),
			("1010101010101010",'0',"101111","0101010101010101"),
			("0101010101010101",'1',"101100","1010101010101010"),
			("0101010101010101",'1',"101100","0101010101010101"),
			("1010101010101010",'1',"101101","0101010101010101"),
			("1010101010101010",'1',"101101","1010101010101010"),
			("1010101010101010",'0',"101000","0101010101010101"),
			("1010101010101010",'0',"101000","0101010101010101"),
			("1010101010101010",'0',"101001","0101010101010101"),
			("1010101010101010",'0',"101010","0101010101010101"),
			("1010101010101010",'0',"101011","0101010101010101"),
			("1010101010101010",'0',"101100","0101010101010101"),
			("1010101010101010",'0',"101101","1010101010101010"),
			("1010101010101010",'0',"101110","0101010101010101"),
			("1010101010101010",'0',"101111","0101010101010101"),
			("0101010101010101",'1',"101101","1010101010101010"),
			("0101010101010101",'1',"101101","0101010101010101"),
			("1010101010101010",'1',"101110","0101010101010101"),
			("1010101010101010",'1',"101110","1010101010101010"),
			("1010101010101010",'0',"101000","0101010101010101"),
			("1010101010101010",'0',"101000","0101010101010101"),
			("1010101010101010",'0',"101001","0101010101010101"),
			("1010101010101010",'0',"101010","0101010101010101"),
			("1010101010101010",'0',"101011","0101010101010101"),
			("1010101010101010",'0',"101100","0101010101010101"),
			("1010101010101010",'0',"101101","0101010101010101"),
			("1010101010101010",'0',"101110","1010101010101010"),
			("1010101010101010",'0',"101111","0101010101010101"),
			("0101010101010101",'1',"101110","1010101010101010"),
			("0101010101010101",'1',"101110","0101010101010101"),
			("1010101010101010",'1',"101111","0101010101010101"),
			("1010101010101010",'1',"101111","1010101010101010"),
			("1010101010101010",'0',"101000","0101010101010101"),
			("1010101010101010",'0',"101000","0101010101010101"),
			("1010101010101010",'0',"101001","0101010101010101"),
			("1010101010101010",'0',"101010","0101010101010101"),
			("1010101010101010",'0',"101011","0101010101010101"),
			("1010101010101010",'0',"101100","0101010101010101"),
			("1010101010101010",'0',"101101","0101010101010101"),
			("1010101010101010",'0',"101110","0101010101010101"),
			("1010101010101010",'0',"101111","1010101010101010"),
			("0101010101010101",'1',"101111","1010101010101010"),
			("0101010101010101",'1',"101111","0101010101010101"),
			("0101010101010101",'0',"101000","0101010101010101"),
			("0101010101010101",'0',"101000","0101010101010101"),
			("0101010101010101",'0',"101001","0101010101010101"),
			("0101010101010101",'0',"101010","0101010101010101"),
			("0101010101010101",'0',"101011","0101010101010101"),
			("0101010101010101",'0',"101100","0101010101010101"),
			("0101010101010101",'0',"101101","0101010101010101"),
			("0101010101010101",'0',"101110","0101010101010101"),
			("0101010101010101",'0',"101111","0101010101010101"),
			("0101010101010101",'0',"000101","0000000000000000"),
			("0101010101010101",'0',"000101","0000000000000000"),
			("0101010101010101",'0',"001101","0000010100100001"),
			("0101010101010101",'0',"010101","0000000000000000"),
			("0101010101010101",'0',"011101","0000000000000000"),
			("0101010101010101",'0',"100101","0000000000000000"),
			("0101010101010101",'0',"101101","0101010101010101"),
			("0101010101010101",'0',"110101","0000000000000000"),
			("0101010101010101",'0',"111101","0000000000000000"),
			("0101010101010101",'1',"000101","0000000000000000"),
			("0101010101010101",'1',"000101","0101010101010101"),
			("0101010101010101",'1',"001101","0000010100100001"),
			("0101010101010101",'1',"001101","0101010101010101"),
			("0101010101010101",'1',"010101","0000000000000000"),
			("0101010101010101",'1',"010101","0101010101010101"),
			("0101010101010101",'1',"011101","0000000000000000"),
			("0101010101010101",'1',"011101","0101010101010101"),
			("0101010101010101",'1',"100101","0000000000000000"),
			("0101010101010101",'1',"100101","0101010101010101"),
			("0101010101010101",'1',"101101","0101010101010101"),
			("0101010101010101",'1',"101101","0101010101010101"),
			("0101010101010101",'1',"110101","0000000000000000"),
			("0101010101010101",'1',"110101","0101010101010101"),
			("0101010101010101",'1',"111101","0000000000000000"),
			("0101010101010101",'1',"111101","0101010101010101"),
			("0101010101010101",'0',"000101","0101010101010101"),
			("0101010101010101",'0',"000101","0101010101010101"),
			("0101010101010101",'0',"001101","0101010101010101"),
			("0101010101010101",'0',"010101","0101010101010101"),
			("0101010101010101",'0',"011101","0101010101010101"),
			("0101010101010101",'0',"100101","0101010101010101"),
			("0101010101010101",'0',"101101","0101010101010101"),
			("0101010101010101",'0',"110101","0101010101010101"),
			("0101010101010101",'0',"111101","0101010101010101"),
			("1010101010101010",'1',"000101","0101010101010101"),
			("1010101010101010",'1',"000101","1010101010101010"),
			("1010101010101010",'0',"000101","1010101010101010"),
			("1010101010101010",'0',"000101","1010101010101010"),
			("1010101010101010",'0',"001101","0101010101010101"),
			("1010101010101010",'0',"010101","0101010101010101"),
			("1010101010101010",'0',"011101","0101010101010101"),
			("1010101010101010",'0',"100101","0101010101010101"),
			("1010101010101010",'0',"101101","0101010101010101"),
			("1010101010101010",'0',"110101","0101010101010101"),
			("1010101010101010",'0',"111101","0101010101010101"),
			("0101010101010101",'1',"000101","1010101010101010"),
			("0101010101010101",'1',"000101","0101010101010101"),
			("1010101010101010",'1',"001101","0101010101010101"),
			("1010101010101010",'1',"001101","1010101010101010"),
			("1010101010101010",'0',"000101","0101010101010101"),
			("1010101010101010",'0',"000101","0101010101010101"),
			("1010101010101010",'0',"001101","1010101010101010"),
			("1010101010101010",'0',"010101","0101010101010101"),
			("1010101010101010",'0',"011101","0101010101010101"),
			("1010101010101010",'0',"100101","0101010101010101"),
			("1010101010101010",'0',"101101","0101010101010101"),
			("1010101010101010",'0',"110101","0101010101010101"),
			("1010101010101010",'0',"111101","0101010101010101"),
			("0101010101010101",'1',"001101","1010101010101010"),
			("0101010101010101",'1',"001101","0101010101010101"),
			("1010101010101010",'1',"010101","0101010101010101"),
			("1010101010101010",'1',"010101","1010101010101010"),
			("1010101010101010",'0',"000101","0101010101010101"),
			("1010101010101010",'0',"000101","0101010101010101"),
			("1010101010101010",'0',"001101","0101010101010101"),
			("1010101010101010",'0',"010101","1010101010101010"),
			("1010101010101010",'0',"011101","0101010101010101"),
			("1010101010101010",'0',"100101","0101010101010101"),
			("1010101010101010",'0',"101101","0101010101010101"),
			("1010101010101010",'0',"110101","0101010101010101"),
			("1010101010101010",'0',"111101","0101010101010101"),
			("0101010101010101",'1',"010101","1010101010101010"),
			("0101010101010101",'1',"010101","0101010101010101"),
			("1010101010101010",'1',"011101","0101010101010101"),
			("1010101010101010",'1',"011101","1010101010101010"),
			("1010101010101010",'0',"000101","0101010101010101"),
			("1010101010101010",'0',"000101","0101010101010101"),
			("1010101010101010",'0',"001101","0101010101010101"),
			("1010101010101010",'0',"010101","0101010101010101"),
			("1010101010101010",'0',"011101","1010101010101010"),
			("1010101010101010",'0',"100101","0101010101010101"),
			("1010101010101010",'0',"101101","0101010101010101"),
			("1010101010101010",'0',"110101","0101010101010101"),
			("1010101010101010",'0',"111101","0101010101010101"),
			("0101010101010101",'1',"011101","1010101010101010"),
			("0101010101010101",'1',"011101","0101010101010101"),
			("1010101010101010",'1',"100101","0101010101010101"),
			("1010101010101010",'1',"100101","1010101010101010"),
			("1010101010101010",'0',"000101","0101010101010101"),
			("1010101010101010",'0',"000101","0101010101010101"),
			("1010101010101010",'0',"001101","0101010101010101"),
			("1010101010101010",'0',"010101","0101010101010101"),
			("1010101010101010",'0',"011101","0101010101010101"),
			("1010101010101010",'0',"100101","1010101010101010"),
			("1010101010101010",'0',"101101","0101010101010101"),
			("1010101010101010",'0',"110101","0101010101010101"),
			("1010101010101010",'0',"111101","0101010101010101"),
			("0101010101010101",'1',"100101","1010101010101010"),
			("0101010101010101",'1',"100101","0101010101010101"),
			("1010101010101010",'1',"101101","0101010101010101"),
			("1010101010101010",'1',"101101","1010101010101010"),
			("1010101010101010",'0',"000101","0101010101010101"),
			("1010101010101010",'0',"000101","0101010101010101"),
			("1010101010101010",'0',"001101","0101010101010101"),
			("1010101010101010",'0',"010101","0101010101010101"),
			("1010101010101010",'0',"011101","0101010101010101"),
			("1010101010101010",'0',"100101","0101010101010101"),
			("1010101010101010",'0',"101101","1010101010101010"),
			("1010101010101010",'0',"110101","0101010101010101"),
			("1010101010101010",'0',"111101","0101010101010101"),
			("0101010101010101",'1',"101101","1010101010101010"),
			("0101010101010101",'1',"101101","0101010101010101"),
			("1010101010101010",'1',"110101","0101010101010101"),
			("1010101010101010",'1',"110101","1010101010101010"),
			("1010101010101010",'0',"000101","0101010101010101"),
			("1010101010101010",'0',"000101","0101010101010101"),
			("1010101010101010",'0',"001101","0101010101010101"),
			("1010101010101010",'0',"010101","0101010101010101"),
			("1010101010101010",'0',"011101","0101010101010101"),
			("1010101010101010",'0',"100101","0101010101010101"),
			("1010101010101010",'0',"101101","0101010101010101"),
			("1010101010101010",'0',"110101","1010101010101010"),
			("1010101010101010",'0',"111101","0101010101010101"),
			("0101010101010101",'1',"110101","1010101010101010"),
			("0101010101010101",'1',"110101","0101010101010101"),
			("1010101010101010",'1',"111101","0101010101010101"),
			("1010101010101010",'1',"111101","1010101010101010"),
			("1010101010101010",'0',"000101","0101010101010101"),
			("1010101010101010",'0',"000101","0101010101010101"),
			("1010101010101010",'0',"001101","0101010101010101"),
			("1010101010101010",'0',"010101","0101010101010101"),
			("1010101010101010",'0',"011101","0101010101010101"),
			("1010101010101010",'0',"100101","0101010101010101"),
			("1010101010101010",'0',"101101","0101010101010101"),
			("1010101010101010",'0',"110101","0101010101010101"),
			("1010101010101010",'0',"111101","1010101010101010"),
			("0101010101010101",'1',"111101","1010101010101010"),
			("0101010101010101",'1',"111101","0101010101010101"),
			("0101010101010101",'0',"000101","0101010101010101"),
			("0101010101010101",'0',"000101","0101010101010101"),
			("0101010101010101",'0',"001101","0101010101010101"),
			("0101010101010101",'0',"010101","0101010101010101"),
			("0101010101010101",'0',"011101","0101010101010101"),
			("0101010101010101",'0',"100101","0101010101010101"),
			("0101010101010101",'0',"101101","0101010101010101"),
			("0101010101010101",'0',"110101","0101010101010101"),
			("0101010101010101",'0',"111101","0101010101010101")
			);
		
	begin

		for i in patterns'range loop
			s_input <= patterns(i).input;
			s_load <= patterns(i).load;
			s_address <= patterns(i).address;
			wait for 40 ns;
			assert s_output = patterns(i).output
			report "bad output" severity error;
		end loop;
	

		assert false report "end of test" severity note;
		s_finished <= '1';	
		wait;
	
	end process;

end architecture RTL;
