library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Ram8_tb is
end entity Ram8_tb;

architecture RTL of Ram8_tb is
	signal s_clk    : std_logic;
	signal s_output : std_logic_vector(15 downto 0);
	signal s_load   : std_logic := '0';
	signal s_input  : std_logic_vector(15 downto 0);
	signal s_finished : std_logic := '0';
	signal s_address : std_logic_vector(2 downto 0);
	
	type pattern_type is record
		input : std_logic_vector(15 downto 0);
		load : std_logic;
		address : std_logic_vector(2 downto 0);
		output : std_logic_vector(15 downto 0);
	end record;
	
	type pattern_array is array (natural range <>) of pattern_type;
	
	
begin
	clock_inst : entity work.ClockGenerator
		generic map(PERIOD => 20 ns)
		port map(finished => s_finished,
		clk => s_clk);

	RAM8: entity work.Ram8
		port map(
			clk     => s_clk,
			rst     => '0',
			load    => s_load,
			address => s_address,
			input   => s_input,
			output  => s_output
		);
	
	process
		constant patterns : pattern_array := (
			("0000000000000000",'0',"000","0000000000000000"),
			("0000000000000000",'0',"000","0000000000000000"),
			("0000000000000000",'1',"000","0000000000000000"),
			("0000000000000000",'1',"000","0000000000000000"),
			("0010101101100111",'0',"000","0000000000000000"),
			("0010101101100111",'0',"000","0000000000000000"),
			("0010101101100111",'1',"001","0000000000000000"),
			("0010101101100111",'1',"001","0010101101100111"),
			("0010101101100111",'0',"000","0000000000000000"),
			("0010101101100111",'0',"000","0000000000000000"),
			("0000110100000101",'0',"011","0000000000000000"),
			("0000110100000101",'0',"011","0000000000000000"),
			("0000110100000101",'1',"011","0000000000000000"),
			("0000110100000101",'1',"011","0000110100000101"),
			("0000110100000101",'0',"011","0000110100000101"),
			("0000110100000101",'0',"011","0000110100000101"),
			("0000110100000101",'0',"001","0010101101100111"),
			("0001111001100001",'0',"001","0010101101100111"),
			("0001111001100001",'0',"001","0010101101100111"),
			("0001111001100001",'1',"111","0000000000000000"),
			("0001111001100001",'1',"111","0001111001100001"),
			("0001111001100001",'0',"111","0001111001100001"),
			("0001111001100001",'0',"111","0001111001100001"),
			("0001111001100001",'0',"011","0000110100000101"),
			("0001111001100001",'0',"111","0001111001100001"),
			("0001111001100001",'0',"000","0000000000000000"),
			("0001111001100001",'0',"000","0000000000000000"),
			("0001111001100001",'0',"001","0010101101100111"),
			("0001111001100001",'0',"010","0000000000000000"),
			("0001111001100001",'0',"011","0000110100000101"),
			("0001111001100001",'0',"100","0000000000000000"),
			("0001111001100001",'0',"101","0000000000000000"),
			("0001111001100001",'0',"110","0000000000000000"),
			("0001111001100001",'0',"111","0001111001100001"),
			("0101010101010101",'1',"000","0000000000000000"),
			("0101010101010101",'1',"000","0101010101010101"),
			("0101010101010101",'1',"001","0010101101100111"),
			("0101010101010101",'1',"001","0101010101010101"),
			("0101010101010101",'1',"010","0000000000000000"),
			("0101010101010101",'1',"010","0101010101010101"),
			("0101010101010101",'1',"011","0000110100000101"),
			("0101010101010101",'1',"011","0101010101010101"),
			("0101010101010101",'1',"100","0000000000000000"),
			("0101010101010101",'1',"100","0101010101010101"),
			("0101010101010101",'1',"101","0000000000000000"),
			("0101010101010101",'1',"101","0101010101010101"),
			("0101010101010101",'1',"110","0000000000000000"),
			("0101010101010101",'1',"110","0101010101010101"),
			("0101010101010101",'1',"111","0001111001100001"),
			("0101010101010101",'1',"111","0101010101010101"),
			("0101010101010101",'0',"000","0101010101010101"),
			("0101010101010101",'0',"000","0101010101010101"),
			("0101010101010101",'0',"001","0101010101010101"),
			("0101010101010101",'0',"010","0101010101010101"),
			("0101010101010101",'0',"011","0101010101010101"),
			("0101010101010101",'0',"100","0101010101010101"),
			("0101010101010101",'0',"101","0101010101010101"),
			("0101010101010101",'0',"110","0101010101010101"),
			("0101010101010101",'0',"111","0101010101010101"),
			("1010101010101010",'1',"000","0101010101010101"),
			("1010101010101010",'1',"000","1010101010101010"),
			("1010101010101010",'0',"000","1010101010101010"),
			("1010101010101010",'0',"000","1010101010101010"),
			("1010101010101010",'0',"001","0101010101010101"),
			("1010101010101010",'0',"010","0101010101010101"),
			("1010101010101010",'0',"011","0101010101010101"),
			("1010101010101010",'0',"100","0101010101010101"),
			("1010101010101010",'0',"101","0101010101010101"),
			("1010101010101010",'0',"110","0101010101010101"),
			("1010101010101010",'0',"111","0101010101010101"),
			("0101010101010101",'1',"000","1010101010101010"),
			("0101010101010101",'1',"000","0101010101010101"),
			("1010101010101010",'1',"001","0101010101010101"),
			("1010101010101010",'1',"001","1010101010101010"),
			("1010101010101010",'0',"000","0101010101010101"),
			("1010101010101010",'0',"000","0101010101010101"),
			("1010101010101010",'0',"001","1010101010101010"),
			("1010101010101010",'0',"010","0101010101010101"),
			("1010101010101010",'0',"011","0101010101010101"),
			("1010101010101010",'0',"100","0101010101010101"),
			("1010101010101010",'0',"101","0101010101010101"),
			("1010101010101010",'0',"110","0101010101010101"),
			("1010101010101010",'0',"111","0101010101010101"),
			("0101010101010101",'1',"001","1010101010101010"),
			("0101010101010101",'1',"001","0101010101010101"),
			("1010101010101010",'1',"010","0101010101010101"),
			("1010101010101010",'1',"010","1010101010101010"),
			("1010101010101010",'0',"000","0101010101010101"),
			("1010101010101010",'0',"000","0101010101010101"),
			("1010101010101010",'0',"001","0101010101010101"),
			("1010101010101010",'0',"010","1010101010101010"),
			("1010101010101010",'0',"011","0101010101010101"),
			("1010101010101010",'0',"100","0101010101010101"),
			("1010101010101010",'0',"101","0101010101010101"),
			("1010101010101010",'0',"110","0101010101010101"),
			("1010101010101010",'0',"111","0101010101010101"),
			("0101010101010101",'1',"010","1010101010101010"),
			("0101010101010101",'1',"010","0101010101010101"),
			("1010101010101010",'1',"011","0101010101010101"),
			("1010101010101010",'1',"011","1010101010101010"),
			("1010101010101010",'0',"000","0101010101010101"),
			("1010101010101010",'0',"000","0101010101010101"),
			("1010101010101010",'0',"001","0101010101010101"),
			("1010101010101010",'0',"010","0101010101010101"),
			("1010101010101010",'0',"011","1010101010101010"),
			("1010101010101010",'0',"100","0101010101010101"),
			("1010101010101010",'0',"101","0101010101010101"),
			("1010101010101010",'0',"110","0101010101010101"),
			("1010101010101010",'0',"111","0101010101010101"),
			("0101010101010101",'1',"011","1010101010101010"),
			("0101010101010101",'1',"011","0101010101010101"),
			("1010101010101010",'1',"100","0101010101010101"),
			("1010101010101010",'1',"100","1010101010101010"),
			("1010101010101010",'0',"000","0101010101010101"),
			("1010101010101010",'0',"000","0101010101010101"),
			("1010101010101010",'0',"001","0101010101010101"),
			("1010101010101010",'0',"010","0101010101010101"),
			("1010101010101010",'0',"011","0101010101010101"),
			("1010101010101010",'0',"100","1010101010101010"),
			("1010101010101010",'0',"101","0101010101010101"),
			("1010101010101010",'0',"110","0101010101010101"),
			("1010101010101010",'0',"111","0101010101010101"),
			("0101010101010101",'1',"100","1010101010101010"),
			("0101010101010101",'1',"100","0101010101010101"),
			("1010101010101010",'1',"101","0101010101010101"),
			("1010101010101010",'1',"101","1010101010101010"),
			("1010101010101010",'0',"000","0101010101010101"),
			("1010101010101010",'0',"000","0101010101010101"),
			("1010101010101010",'0',"001","0101010101010101"),
			("1010101010101010",'0',"010","0101010101010101"),
			("1010101010101010",'0',"011","0101010101010101"),
			("1010101010101010",'0',"100","0101010101010101"),
			("1010101010101010",'0',"101","1010101010101010"),
			("1010101010101010",'0',"110","0101010101010101"),
			("1010101010101010",'0',"111","0101010101010101"),
			("0101010101010101",'1',"101","1010101010101010"),
			("0101010101010101",'1',"101","0101010101010101"),
			("1010101010101010",'1',"110","0101010101010101"),
			("1010101010101010",'1',"110","1010101010101010"),
			("1010101010101010",'0',"000","0101010101010101"),
			("1010101010101010",'0',"000","0101010101010101"),
			("1010101010101010",'0',"001","0101010101010101"),
			("1010101010101010",'0',"010","0101010101010101"),
			("1010101010101010",'0',"011","0101010101010101"),
			("1010101010101010",'0',"100","0101010101010101"),
			("1010101010101010",'0',"101","0101010101010101"),
			("1010101010101010",'0',"110","1010101010101010"),
			("1010101010101010",'0',"111","0101010101010101"),
			("0101010101010101",'1',"110","1010101010101010"),
			("0101010101010101",'1',"110","0101010101010101"),
			("1010101010101010",'1',"111","0101010101010101"),
			("1010101010101010",'1',"111","1010101010101010"),
			("1010101010101010",'0',"000","0101010101010101"),
			("1010101010101010",'0',"000","0101010101010101"),
			("1010101010101010",'0',"001","0101010101010101"),
			("1010101010101010",'0',"010","0101010101010101"),
			("1010101010101010",'0',"011","0101010101010101"),
			("1010101010101010",'0',"100","0101010101010101"),
			("1010101010101010",'0',"101","0101010101010101"),
			("1010101010101010",'0',"110","0101010101010101"),
			("1010101010101010",'0',"111","1010101010101010"),
			("0101010101010101",'1',"111","1010101010101010"),
			("0101010101010101",'1',"111","0101010101010101"),
			("0101010101010101",'0',"000","0101010101010101"),
			("0101010101010101",'0',"000","0101010101010101"),
			("0101010101010101",'0',"001","0101010101010101"),
			("0101010101010101",'0',"010","0101010101010101"),
			("0101010101010101",'0',"011","0101010101010101"),
			("0101010101010101",'0',"100","0101010101010101"),
			("0101010101010101",'0',"101","0101010101010101"),
			("0101010101010101",'0',"110","0101010101010101"),
			("0101010101010101",'0',"111","0101010101010101")
			);
		
	begin

		for i in patterns'range loop
			s_input <= patterns(i).input;
			s_load <= patterns(i).load;
			s_address <= patterns(i).address;
			wait for 20 ns;
			assert s_output = patterns(i).output
			report "bad output" severity error;
		end loop;
	

		assert false report "end of test" severity note;
		s_finished <= '1';	
		wait;
	
	end process;

end architecture RTL;
