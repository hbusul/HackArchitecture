--  A testbench has no ports.
entity Mux4Way16_tb is
end Mux4Way16_tb;

library ieee;
use ieee.std_logic_1164.all;
architecture behav of Mux4Way16_tb is
	type pattern_type is record
		input0 : std_logic_vector(15 downto 0);
		input1 : std_logic_vector(15 downto 0);
		input2 : std_logic_vector(15 downto 0);
		input3 : std_logic_vector(15 downto 0);
		sel    : std_logic_vector(1 downto 0);
		output : std_logic_vector(15 downto 0);
	end record;

	type pattern_array is array (natural range <>) of pattern_type;
	
	component Mux4Way16
		port(
			input0 : in  std_logic_vector(15 downto 0);
			input1 : in  std_logic_vector(15 downto 0);
			input2 : in  std_logic_vector(15 downto 0);
			input3 : in  std_logic_vector(15 downto 0);
			sel    : in  std_logic_vector(1 downto 0);
			output : out std_logic_vector(15 downto 0)
		);
	end component Mux4Way16;


	signal s_input0 : std_logic_vector(15 downto 0);
	signal s_input1 : std_logic_vector(15 downto 0);
	signal s_input2 : std_logic_vector(15 downto 0);
	signal s_input3 : std_logic_vector(15 downto 0);
	signal s_sel    : std_logic_vector(1 downto 0);
	signal s_output : std_logic_vector(15 downto 0);

begin
	
	mux0: Mux4Way16
		port map(
			input0 => s_input0,
			input1 => s_input1,
			input2 => s_input2,
			input3 => s_input3,
			sel    => s_sel,
			output => s_output
		);
	
	process
		constant patterns : pattern_array := (
			("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000",
			"00", "0000000000000000"
			),
			("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000",
			"01", "0000000000000000"
			),
			("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000",
			"10", "0000000000000000"
			),
			("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000",
			"11", "0000000000000000"
			),
			
			("1111111111111111", "1111111111111111", "1111111111111111", "1111111111111111",
			"00", "1111111111111111"
			),
			("1111111111111111", "1111111111111111", "1111111111111111", "1111111111111111",
			"01", "1111111111111111"
			),
			("1111111111111111", "1111111111111111", "1111111111111111", "1111111111111111",
			"10", "1111111111111111"
			),
			("1111111111111111", "1111111111111111", "1111111111111111", "1111111111111111",
			"11", "1111111111111111"
			),
			
			
			("0000000000000000", "1111111111111111", "0000000000000000", "1111111111111111",
			"00", "0000000000000000"
			),
			("0000000000000000", "1111111111111111", "0000000000000000", "1111111111111111",
			"01", "1111111111111111"
			),
			("0000000000000000", "1111111111111111", "0000000000000000", "1111111111111111",
			"10", "0000000000000000"
			),
			("0000000000000000", "1111111111111111", "0000000000000000", "1111111111111111",
			"11", "1111111111111111"
			),
			
			
			("1111111111111111", "0000000000000000", "1111111111111111", "0000000000000000",
			"00", "1111111111111111"
			),
			("1111111111111111", "0000000000000000", "1111111111111111", "0000000000000000",
			"01", "0000000000000000"
			),
			("1111111111111111", "0000000000000000", "1111111111111111", "0000000000000000",
			"10", "1111111111111111"
			),
			("1111111111111111", "0000000000000000", "1111111111111111", "0000000000000000",
			"11", "0000000000000000"
			),
			
			
			("1010101010110111", "0000000000000000", "1111111111111111", "1101001010101010",
			"00", "1010101010110111"
			),
			("1010101010110111", "0000000000000000", "1111111111111111", "1101001010101010",
			"01", "0000000000000000"
			),
			("1010101010110111", "0000000000000000", "1111111111111111", "1101001010101010",
			"10", "1111111111111111"
			),
			("1010101010110111", "0000000000000000", "1111111111111111", "1101001010101010",
			"11", "1101001010101010"
			),
			
			("0000000000001111", "0000000011110000", "0000111100000000", "1111000000000000",
			"00", "0000000000001111"
			),
			("0000000000001111", "0000000011110000", "0000111100000000", "1111000000000000",
			"01", "0000000011110000"
			),
			("0000000000001111", "0000000011110000", "0000111100000000", "1111000000000000",
			"10", "0000111100000000"
			),
			("0000000000001111", "0000000011110000", "0000111100000000", "1111000000000000",
			"11", "1111000000000000"
			)
		
		);

	begin
		for i in patterns'range loop
			s_input0 <= patterns(i).input0;
			s_input1 <= patterns(i).input1;
			s_input2 <= patterns(i).input2;
			s_input3 <= patterns(i).input3;
			s_sel    <= patterns(i).sel;
			wait for 1 ns;
			assert s_output = patterns(i).output
			report "bad output" severity error;
		end loop;
		assert false report "end of test" severity note;
		wait;
	end process;
end behav;
