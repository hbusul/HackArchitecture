--  A testbench has no ports.
entity Mux8Way16_tb is
end Mux8Way16_tb;

library ieee;
use ieee.std_logic_1164.all;
architecture behav of Mux8Way16_tb is
	type pattern_type is record
		input0 : std_logic_vector(15 downto 0);
		input1 : std_logic_vector(15 downto 0);
		input2 : std_logic_vector(15 downto 0);
		input3 : std_logic_vector(15 downto 0);
		input4 : std_logic_vector(15 downto 0);
		input5 : std_logic_vector(15 downto 0);
		input6 : std_logic_vector(15 downto 0);
		input7 : std_logic_vector(15 downto 0);
		sel    : std_logic_vector(2 downto 0);
		output : std_logic_vector(15 downto 0);
	end record;

	type pattern_array is array (natural range <>) of pattern_type;

	component Mux8Way16
		port(
			input0 : in  std_logic_vector(15 downto 0);
			input1 : in  std_logic_vector(15 downto 0);
			input2 : in  std_logic_vector(15 downto 0);
			input3 : in  std_logic_vector(15 downto 0);
			input4 : in  std_logic_vector(15 downto 0);
			input5 : in  std_logic_vector(15 downto 0);
			input6 : in  std_logic_vector(15 downto 0);
			input7 : in  std_logic_vector(15 downto 0);
			sel    : in  std_logic_vector(2 downto 0);
			output : out std_logic_vector(15 downto 0)
		);
	end component Mux8Way16;

	signal s_input0 : std_logic_vector(15 downto 0);
	signal s_input1 : std_logic_vector(15 downto 0);
	signal s_input2 : std_logic_vector(15 downto 0);
	signal s_input3 : std_logic_vector(15 downto 0);
	signal s_input4 : std_logic_vector(15 downto 0);
	signal s_input5 : std_logic_vector(15 downto 0);
	signal s_input6 : std_logic_vector(15 downto 0);
	signal s_input7 : std_logic_vector(15 downto 0);
	signal s_sel    : std_logic_vector(2 downto 0);
	signal s_output : std_logic_vector(15 downto 0);

begin

	mux0 : component Mux8Way16
		port map(
			input0 => s_input0,
			input1 => s_input1,
			input2 => s_input2,
			input3 => s_input3,
			input4 => s_input4,
			input5 => s_input5,
			input6 => s_input6,
			input7 => s_input7,
			sel    => s_sel,
			output => s_output
		);

	process
		constant patterns : pattern_array := (
			("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000",
		     "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000",	
			 "000", "0000000000000000"),
			("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000",
			 "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000",	
			 "001", "0000000000000000"),
			("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000",
			 "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000",	
			 "010", "0000000000000000"),
			("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000",
			 "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000",	
			 "011", "0000000000000000"),
			("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000",
			 "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000",	
			 "100", "0000000000000000"),
			("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000",
			 "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000",	
			 "101", "0000000000000000"),
			("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000",
			 "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000",	
			 "110", "0000000000000000"),
			("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000",
			 "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000",	
			 "111", "0000000000000000"),
			 
			
			("1111111111111111", "1111111111111111", "1111111111111111", "1111111111111111",
			 "1111111111111111", "1111111111111111", "1111111111111111", "1111111111111111",	
			 "000", "1111111111111111"),
			("1111111111111111", "1111111111111111", "1111111111111111", "1111111111111111",
			 "1111111111111111", "1111111111111111", "1111111111111111", "1111111111111111",	
			 "001", "1111111111111111"),
			("1111111111111111", "1111111111111111", "1111111111111111", "1111111111111111",
			 "1111111111111111", "1111111111111111", "1111111111111111", "1111111111111111",	
			 "010", "1111111111111111"),
			("1111111111111111", "1111111111111111", "1111111111111111", "1111111111111111",
			 "1111111111111111", "1111111111111111", "1111111111111111", "1111111111111111",	
			 "011", "1111111111111111"),
			("1111111111111111", "1111111111111111", "1111111111111111", "1111111111111111",
			 "1111111111111111", "1111111111111111", "1111111111111111", "1111111111111111",	
			 "100", "1111111111111111"),
			("1111111111111111", "1111111111111111", "1111111111111111", "1111111111111111",
			 "1111111111111111", "1111111111111111", "1111111111111111", "1111111111111111",	
			 "101", "1111111111111111"),
			("1111111111111111", "1111111111111111", "1111111111111111", "1111111111111111",
			 "1111111111111111", "1111111111111111", "1111111111111111", "1111111111111111",	
			 "110", "1111111111111111"),
			("1111111111111111", "1111111111111111", "1111111111111111", "1111111111111111",
			 "1111111111111111", "1111111111111111", "1111111111111111", "1111111111111111",	
			 "111", "1111111111111111"),
			 
			
			("0000000000000000", "1111111111111111", "0000000000000000", "1111111111111111",
			 "0000000000000000", "1111111111111111", "0000000000000000", "1111111111111111",
			 "000", "0000000000000000"),
			("0000000000000000", "1111111111111111", "0000000000000000", "1111111111111111",
			 "0000000000000000", "1111111111111111", "0000000000000000", "1111111111111111",
			 "001", "1111111111111111"),
			("0000000000000000", "1111111111111111", "0000000000000000", "1111111111111111",
			 "0000000000000000", "1111111111111111", "0000000000000000", "1111111111111111",
			 "010", "0000000000000000"),
			("0000000000000000", "1111111111111111", "0000000000000000", "1111111111111111",
			 "0000000000000000", "1111111111111111", "0000000000000000", "1111111111111111",
			 "011", "1111111111111111"),
			("0000000000000000", "1111111111111111", "0000000000000000", "1111111111111111",
			 "0000000000000000", "1111111111111111", "0000000000000000", "1111111111111111",
			 "100", "0000000000000000"),
			("0000000000000000", "1111111111111111", "0000000000000000", "1111111111111111",
			 "0000000000000000", "1111111111111111", "0000000000000000", "1111111111111111",
			 "101", "1111111111111111"),
			("0000000000000000", "1111111111111111", "0000000000000000", "1111111111111111",
			 "0000000000000000", "1111111111111111", "0000000000000000", "1111111111111111",
			 "110", "0000000000000000"),
			("0000000000000000", "1111111111111111", "0000000000000000", "1111111111111111",
			 "0000000000000000", "1111111111111111", "0000000000000000", "1111111111111111",
			 "111", "1111111111111111"),
			  					                     
			 ("1010101010110111", "0000011100100000", "1111111111111111", "1101001010101010",
			  "1010111110110111", "0100001111100000", "0000000000000000", "0001001010100010",
			  "000", "1010101010110111"),
			 ("1010101010110111", "0000011100100000", "1111111111111111", "1101001010101010",
			  "1010111110110111", "0100001111100000", "0000000000000000", "0001001010100010",
			  "001", "0000011100100000"),
			 ("1010101010110111", "0000011100100000", "1111111111111111", "1101001010101010",
			  "1010111110110111", "0100001111100000", "0000000000000000", "0001001010100010",
			  "010", "1111111111111111"),
			 ("1010101010110111", "0000011100100000", "1111111111111111", "1101001010101010",
			  "1010111110110111", "0100001111100000", "0000000000000000", "0001001010100010",
			  "011", "1101001010101010"),
			 ("1010101010110111", "0000011100100000", "1111111111111111", "1101001010101010",
			  "1010111110110111", "0100001111100000", "0000000000000000", "0001001010100010",
			  "100", "1010111110110111"),
			 ("1010101010110111", "0000011100100000", "1111111111111111", "1101001010101010",
			  "1010111110110111", "0100001111100000", "0000000000000000", "0001001010100010",
			  "101", "0100001111100000"),
			 ("1010101010110111", "0000011100100000", "1111111111111111", "1101001010101010",
			  "1010111110110111", "0100001111100000", "0000000000000000", "0001001010100010",
			  "110", "0000000000000000"),
			 ("1010101010110111", "0000011100100000", "1111111111111111", "1101001010101010",
			  "1010111110110111", "0100001111100000", "0000000000000000", "0001001010100010",
			  "111", "0001001010100010")  
			
		);

	begin
		for i in patterns'range loop
			s_input0 <= patterns(i).input0;
			s_input1 <= patterns(i).input1;
			s_input2 <= patterns(i).input2;
			s_input3 <= patterns(i).input3;
			s_input4 <= patterns(i).input4;
			s_input5 <= patterns(i).input5;
			s_input6 <= patterns(i).input6;
			s_input7 <= patterns(i).input7;
			s_sel    <= patterns(i).sel;
			wait for 1 ns;
			assert s_output = patterns(i).output
			report "bad output" severity error;
		end loop;
		assert false report "end of test" severity note;
		wait;
	end process;
end behav;
