library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ALU_tb is
end entity ALU_tb;

architecture behav of ALU_tb is
	signal s_x, s_y                          : std_logic_vector(15 downto 0);
	signal s_zx, s_nx, s_zy, s_ny, s_f, s_no : std_logic;
	signal s_output                          : std_logic_vector(15 downto 0);
	signal s_zr, s_ng                        : std_logic;

	type pattern_type is record
		x, y                  : std_logic_vector(15 downto 0);
		zx, nx, zy, ny, f, no : std_logic;
		output                : std_logic_vector(15 downto 0);
		zr, ng                : std_logic;
	end record;

	type pattern_array is array (natural range <>) of pattern_type;

	component ALU
		port(
			x                     : in  std_logic_vector(15 downto 0);
			y                     : in  std_logic_vector(15 downto 0);
			zx, nx, zy, ny, f, no : in  std_logic;
			output                : out std_logic_vector(15 downto 0);
			zr                    : out std_logic;
			ng                    : out std_logic
		);
	end component ALU;

begin
	alu0 : component ALU
		port map(
			x      => s_x,
			y      => s_y,
			zx     => s_zx,
			nx     => s_nx,
			zy     => s_zy,
			ny     => s_ny,
			f      => s_f,
			no     => s_no,
			output => s_output,
			zr     => s_zr,
			ng     => s_ng
		);

	process
		constant patterns : pattern_array := (
			("0000000000000000", "1111111111111111", '1', '0', '1', '0', '1', '0', "0000000000000000", '1', '0'),
			("0000000000000000", "1111111111111111", '1', '1', '1', '1', '1', '1', "0000000000000001", '0', '0'),
			("0000000000000000", "1111111111111111", '1', '1', '1', '0', '1', '0', "1111111111111111", '0', '1'),
			("0000000000000000", "1111111111111111", '0', '0', '1', '1', '0', '0', "0000000000000000", '1', '0'),
			("0000000000000000", "1111111111111111", '1', '1', '0', '0', '0', '0', "1111111111111111", '0', '1'),
			("0000000000000000", "1111111111111111", '0', '0', '1', '1', '0', '1', "1111111111111111", '0', '1'),
			("0000000000000000", "1111111111111111", '1', '1', '0', '0', '0', '1', "0000000000000000", '1', '0'),
			("0000000000000000", "1111111111111111", '0', '0', '1', '1', '1', '1', "0000000000000000", '1', '0'),
			("0000000000000000", "1111111111111111", '1', '1', '0', '0', '1', '1', "0000000000000001", '0', '0'),
			("0000000000000000", "1111111111111111", '0', '1', '1', '1', '1', '1', "0000000000000001", '0', '0'),
			("0000000000000000", "1111111111111111", '1', '1', '0', '1', '1', '1', "0000000000000000", '1', '0'),
			("0000000000000000", "1111111111111111", '0', '0', '1', '1', '1', '0', "1111111111111111", '0', '1'),
			("0000000000000000", "1111111111111111", '1', '1', '0', '0', '1', '0', "1111111111111110", '0', '1'),
			("0000000000000000", "1111111111111111", '0', '0', '0', '0', '1', '0', "1111111111111111", '0', '1'),
			("0000000000000000", "1111111111111111", '0', '1', '0', '0', '1', '1', "0000000000000001", '0', '0'),
			("0000000000000000", "1111111111111111", '0', '0', '0', '1', '1', '1', "1111111111111111", '0', '1'),
			("0000000000000000", "1111111111111111", '0', '0', '0', '0', '0', '0', "0000000000000000", '1', '0'),
			("0000000000000000", "1111111111111111", '0', '1', '0', '1', '0', '1', "1111111111111111", '0', '1'),
			("0000000000010001", "0000000000000011", '1', '0', '1', '0', '1', '0', "0000000000000000", '1', '0'),
			("0000000000010001", "0000000000000011", '1', '1', '1', '1', '1', '1', "0000000000000001", '0', '0'),
			("0000000000010001", "0000000000000011", '1', '1', '1', '0', '1', '0', "1111111111111111", '0', '1'),
			("0000000000010001", "0000000000000011", '0', '0', '1', '1', '0', '0', "0000000000010001", '0', '0'),
			("0000000000010001", "0000000000000011", '1', '1', '0', '0', '0', '0', "0000000000000011", '0', '0'),
			("0000000000010001", "0000000000000011", '0', '0', '1', '1', '0', '1', "1111111111101110", '0', '1'),
			("0000000000010001", "0000000000000011", '1', '1', '0', '0', '0', '1', "1111111111111100", '0', '1'),
			("0000000000010001", "0000000000000011", '0', '0', '1', '1', '1', '1', "1111111111101111", '0', '1'),
			("0000000000010001", "0000000000000011", '1', '1', '0', '0', '1', '1', "1111111111111101", '0', '1'),
			("0000000000010001", "0000000000000011", '0', '1', '1', '1', '1', '1', "0000000000010010", '0', '0'),
			("0000000000010001", "0000000000000011", '1', '1', '0', '1', '1', '1', "0000000000000100", '0', '0'),
			("0000000000010001", "0000000000000011", '0', '0', '1', '1', '1', '0', "0000000000010000", '0', '0'),
			("0000000000010001", "0000000000000011", '1', '1', '0', '0', '1', '0', "0000000000000010", '0', '0'),
			("0000000000010001", "0000000000000011", '0', '0', '0', '0', '1', '0', "0000000000010100", '0', '0'),
			("0000000000010001", "0000000000000011", '0', '1', '0', '0', '1', '1', "0000000000001110", '0', '0'),
			("0000000000010001", "0000000000000011", '0', '0', '0', '1', '1', '1', "1111111111110010", '0', '1'),
			("0000000000010001", "0000000000000011", '0', '0', '0', '0', '0', '0', "0000000000000001", '0', '0'),
			("0000000000010001", "0000000000000011", '0', '1', '0', '1', '0', '1', "0000000000010011", '0', '0')
		);
	begin
		for i in patterns'range loop
			s_x <= patterns(i).x;
			s_y <= patterns(i).y;
			s_zx <= patterns(i).zx;
			s_nx <= patterns(i).nx;
			s_zy <= patterns(i).zy;
			s_ny <= patterns(i).ny;
			s_f <= patterns(i).f;
			s_no <= patterns(i).no;
			
			wait for 1 ns;
			assert s_output = patterns(i).output
			report "bad output" severity error;
			
			assert s_zr = patterns(i).zr
			report "bad zr" severity error;
			
			assert s_ng = patterns(i).ng
			report "bad ng" severity error;
		end loop;
		
		assert false report "end of test" severity note;
		wait;
		
	end process;

end architecture behav;
